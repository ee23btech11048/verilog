module universal_shift_reg (
    input clk,
    input rst_n,
    input [8:0] select,
    input [15:0] parallel_in,
    input serial_left_data_in,
    input serial_right_data_in,
    output reg [15:0] p_dout,
    output s_left_dout,
    output s_right_dout
);

// Define parameters, instantiate shift register modules, and define default behavior

endmodule

